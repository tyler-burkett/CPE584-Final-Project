{?header?}

`celldefine
`timescale {?timescale?}


module {?lib?}_a221o_{?drive?}  (
output {?in0?},

input {?in0?},
input {?in1?},
input {?in2?},
input {?in3?},
input {?in4?}

`ifdef SC_USE_PG_PIN
, input {?vpwr0?}
, input {?vgnd0?}
, input {?vpb0?}
, input {?vnb0?}
`endif

);

`ifdef functional
`else
`ifdef SC_USE_PG_PIN
`else
supply1 {?vpwr0?};
supply0 {?vgnd0?};
supply1 {?vpb0?};
supply0 {?vnb0?};
`endif
`endif


  wire csi_opt_273;
  wire csi_opt_274;

`ifdef functional
`else
reg csi_notifier;

	specify
		({?in0?} +=> {?in0?}) =  (0:0:0,0:0:0);
		({?in0?} -=> {?in0?}) =  (0:0:0,0:0:0);
		({?in1?} +=> {?in0?}) =  (0:0:0,0:0:0);
		({?in1?} -=> {?in0?}) =  (0:0:0,0:0:0);
		({?in2?} +=> {?in0?}) =  (0:0:0,0:0:0);
		({?in2?} -=> {?in0?}) =  (0:0:0,0:0:0);
		({?in3?} +=> {?in0?}) =  (0:0:0,0:0:0);
		({?in3?} -=> {?in0?}) =  (0:0:0,0:0:0);
		({?in4?} +=> {?in0?}) =  (0:0:0,0:0:0);
		({?in4?} -=> {?in0?}) =  (0:0:0,0:0:0);
	endspecify
`endif

  and ( csi_opt_273 , {?in2?} , {?in3?} ) ;
  and ( csi_opt_274 , {?in0?} , {?in1?} ) ;
  or  ( UDP_IN_X , csi_opt_274 , csi_opt_273 , {?in4?} ) ;
  `ifdef SC_USE_PG_PIN

  {?lib?}_pg_U_VPWR_VGND (UDP_OUT_X, UDP_IN_X, {?vpwr0?}, {?vgnd0?}) ;
  buf  ({?in0?}, UDP_OUT_X) ;
  `else
    buf ( {?in0?} , UDP_IN_X ) ;
  `endif
endmodule
`endcelldefine
