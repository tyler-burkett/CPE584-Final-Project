{#
	DESCRIPTION
		One 2-input and & one inverted input into 2-input nor
	PARAMETER MAPPING
		in[0]	:	A1
		in[1]	:	A2
		in[2]	:	B1N
		out[0]	:	Y
-#}


{? header ?}


`celldefine
`timescale 1ns / 1ps


module {? lib ?}_{? name ?}_{? drive ?}  (
output {? out[0] ?},

input {? in[0] ?},
input {? in[1] ?},
input {? in[2] ?}

`ifdef SC_USE_PG_PIN
, input {? vpwr[0] ?}
, input {? vgnd[0] ?}
, input {? vpb[0] ?}
, input {? vnb[0] ?}
`endif

);

`ifdef functional
`else
`ifdef SC_USE_PG_PIN
`else
supply1 {? vpwr[0] ?};
supply0 {? vgnd[0] ?};
supply1 {? vpb[0] ?};
supply0 {? vnb[0] ?};
`endif
`endif

  wire b;
   not (b,{? in[2] ?});
   and ( csi_opt_273 , {? in[0] ?} , {? in[1] ?} ) ;
   nor  ( UDP_IN_Y , b , csi_opt_273 ) ;
  `ifdef SC_USE_PG_PIN

  {? lib ?}_pg_U_VPWR_VGND (UDP_OUT_Y, UDP_IN_Y, {? vpwr[0] ?}, {? vgnd[0] ?}) ;
  buf  ({? out[0] ?}, UDP_OUT_Y) ;
  `else
    buf ( {? out[0] ?} , UDP_IN_Y ) ;
  `endif
// modification by B1NB, based on SPR13943.  need to have
`ifdef functional
`else
reg csi_notifier;

        specify
		({? in[0] ?} +=> {? out[0] ?}) =   (0:0:0,0:0:0);
		({? in[0] ?} -=> {? out[0] ?}) =   (0:0:0,0:0:0);
		({? in[1] ?} +=> {? out[0] ?}) =   (0:0:0,0:0:0);
		({? in[1] ?} -=> {? out[0] ?}) =   (0:0:0,0:0:0);
		({? in[2] ?} +=> {? out[0] ?}) =   (0:0:0,0:0:0);
		({? in[2] ?} -=> {? out[0] ?}) =   (0:0:0,0:0:0);
	endspecify
`endif
   
endmodule
`endcelldefine
