{?header?}

`celldefine
`timescale {?timescale?}



module {?lib?}_decap_{?drive?}  (

`ifdef SC_USE_PG_PIN
input {?vpwr0?},
input {?vgnd0?},
input {?vpb0?},
input {?vnb0?}
`endif

);

`ifdef functional
`else
`ifdef SC_USE_PG_PIN
`else
supply1 {?vpwr0?};
supply0 {?vgnd0?};
supply1 {?vpb0?};
supply0 {?vnb0?};
`endif
`endif


endmodule
`endcelldefine
